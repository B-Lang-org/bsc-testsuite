package Bits where

import Vector
import BuildVector

class MyBits a n | a -> n where
  mypack   :: a -> Bit n
  myunpack :: Bit n -> a

instance MyBits (Bit n) n where
  mypack = id
  myunpack = id

instance (Generic a r, MyBits' r n) => MyBits a n where
  mypack   x  = mypack' $ from x
  myunpack bs = to $ myunpack' bs

class MyBits' r n | r -> n where
  mypack'   :: r -> Bit n
  myunpack' :: Bit n -> r

instance (Log ncons ntag, ConBits r ndata, Add ntag ndata n) =>
         MyBits' (MetaData name pkg ncons r) n where
  mypack' (MetaData x) =
    let (tagNum, dat) = packCon x
        tag = pack ((fromInteger tagNum) :: UInt ntag)
    in tag ++ dat
  myunpack' bs =
    let (tag, dat) = split bs
    in MetaData $ unpackCon (primUIntBitsToInteger (tag :: Bit ntag)) dat

class ConBits r n | r -> n where
  packCon   :: r -> (Integer, Bit n)
  unpackCon :: Integer -> Bit n -> r

instance (ConBits a1 n1, ConBits a2 n2, Max n1 n2 n, Add p1 n1 n, Add p2 n2 n) =>
         ConBits (Either a1 a2) n where
  packCon (Left x) =
    let (tag, bs) = packCon x
    in (tag, extend bs)
  packCon (Right x) =
    let (tag, bs) = packCon x
    in (tag, extend bs)
  unpackCon 0 bs = Left $ unpackCon 0 (truncate bs)
  unpackCon i bs = Right $ unpackCon (i - 1) (truncate bs)

instance (MyBits' r n) => ConBits (MetaConsNamed name idx nfields r) n where
  packCon (MetaConsNamed x) = (valueOf idx, mypack' x)
  unpackCon _ bs = MetaConsNamed $ myunpack' bs

instance (MyBits' r n) => ConBits (MetaConsAnon name idx nfields r) n where
  packCon (MetaConsAnon x) = (valueOf idx, mypack' x)
  unpackCon _ bs = MetaConsAnon $ myunpack' bs

instance (MyBits' r1 n1, MyBits' r2 n2, Add n1 n2 n) => MyBits' (r1, r2) n where
  mypack' (x, y) = mypack' x ++ mypack' y
  myunpack' bs = let (bs1, bs2) = split bs
                 in (myunpack' bs1, myunpack' bs2)

instance  MyBits' () 0 where
  mypack' () = 0'b0
  myunpack' _ = ()

instance (MyBits' r n) => MyBits' (MetaField name idx r) n where
  mypack' (MetaField x) = mypack' x
  myunpack' bs = MetaField $ myunpack' bs

instance (MyBits' a m, Bits (Vector n (Bit m)) l) =>
         MyBits' (MetaData name pkg 1 (Vector n a)) l where
  mypack' (MetaData v) = pack $ map mypack' v
  myunpack' = MetaData `compose` map myunpack' `compose` unpack

instance (MyBits a n) => MyBits' (Conc a) n where
  mypack' (Conc x) = mypack x
  myunpack' bs = Conc $ myunpack bs

data Foo = A (UInt 8)
         | B (UInt 16) Bool Bar
         | C
  deriving (Generic, FShow)

struct Bar =
  x :: (UInt 8)
  y :: (UInt 8)
 deriving (Generic, FShow)


data MyUInt n = UInt (Bit n)
  deriving (Generic)

foo :: Vector 3 Foo
foo = vec (A 5) (B 1223 True (Bar {x=42; y=54})) C

fooPack :: Bit 105
fooPack = mypack foo

fooUnpack :: Vector 3 Foo
fooUnpack = myunpack fooPack

sysBits :: Module Empty
sysBits = module
  rules
    when True ==> do
      $display (fshow foo)
      -- $display (fshow fooPack)
      $display (fshow fooUnpack)
      $finish
