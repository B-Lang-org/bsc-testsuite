package GenericTests where

import ListN
import Vector
import BuildVector

-- Represents "evidence" for type equality between a and b,
-- can only be constructed by refl ("reflexive") when a and b are equal.
-- This could move to a library, I suppose?
data TypeEq a b = Refl__
refl :: TypeEq a a
refl = Refl__


data Foo = A (UInt 8) Bool Bar
         | B (UInt 16)
         | C
         | D {a :: (UInt 8); b :: Foo}
  deriving (Eq, FShow)

struct Bar =
  foo :: Foo
  x :: (UInt 8)
 deriving (Eq, FShow)

data Baz a = Baz a a
  deriving (Eq, FShow)

-- Test generic representations
fooRepr :: (Generic Foo r) => TypeEq r
  (Meta (MetaData "Foo" "GenericTests" 4)
   (Either
    (Meta (MetaConsAnon "A" 0 3)
     (Meta (MetaField "_0" 0) (Conc (UInt 8)),
      Meta (MetaField "_1" 1) (Conc Bool),
      Meta (MetaField "_2" 2) (Conc Bar)))
    (Either
     (Meta (MetaConsAnon "B" 1 1)
      (Meta (MetaField "_0" 0) (Conc (UInt 16))))
     (Either (Meta (MetaConsAnon "C" 2 0) ())
      (Meta (MetaConsNamed "D" 3 2)
       (Meta (MetaField "a" 0) (Conc (UInt 8)),
        Meta (MetaField "b" 1) (Conc Foo)))))))
fooRepr = refl

barRepr :: (Generic Bar r) => TypeEq r
  (Meta (MetaData "Bar" "GenericTests" 1)
   (Meta (MetaConsNamed "Bar" 0 2)
    (Meta (MetaField "foo" 0) (Conc Foo),
     Meta (MetaField "x" 1) (Conc (UInt 8)))))
barRepr = refl

bazRepr :: (Generic (Baz a) r) => TypeEq r
  (Meta (MetaData "Baz" "GenericTests" 1)
   (Meta (MetaConsAnon "Baz" 0 2)
    (Meta (MetaField "_0" 0) (Conc a),
     Meta (MetaField "_1" 1) (Conc a))))
bazRepr = refl

bazFooRepr :: (Generic (Baz Foo) r) => TypeEq r
  (Meta (MetaData "Baz" "GenericTests" 1)
   (Meta (MetaConsAnon "Baz" 0 2)
    (Meta (MetaField "_0" 0) (Conc Foo),
     Meta (MetaField "_1" 1) (Conc Foo))))
bazFooRepr = refl

barVec3Repr :: (Generic (Vector 3 Bar) r) => TypeEq r
  (Meta (MetaData "Vector" "Vector" 1) (Vector 3 (Conc Bar)))
barVec3Repr = refl

barListN3Repr :: (Generic (ListN 3 Bar) r) => TypeEq r
  (Meta (MetaData "ListN" "ListN" 1) (Vector 3 (Conc Bar)))
barListN3Repr = refl

-- Test to/from
actTestGeneric :: (Generic a r, FShow a, FShow r, Eq a) => a -> Action
actTestGeneric x = do
  $display "Representation for " (fshow x)
  $display (fshow (from x))
  let res :: a = to (from x)
  if res == x
    then $display "from matches"
    else $display "from mismatch: " (fshow res)

sysGenericTests :: Module Empty
sysGenericTests = module
  rules
    when True ==> do
      actTestGeneric (42 :: UInt 8)
      actTestGeneric (Bar {x=42; foo=C})
      actTestGeneric (A 12 True (Bar {foo=D {a=34; b=C}; x=42}))
      actTestGeneric (Baz C (A 12 True (Bar {foo=D {a=34; b=C}; x=42})))
      actTestGeneric ((vec (Bar {x=42; foo=C}) (Bar {x=3; foo=B 2323})) :: Vector 2 Bar)
--    actTestGeneric ((Bar {x=42; foo=C}) :> (Bar {x=3; foo=B 2323}) :> ListN.nil) -- XXX ListN doesn't have FShow
      $finish
