package UndefinedAttrib where

a :: Attributes__
a = _

m :: Module Empty
m = module
  interface

sysUndefinedAttrib :: Module Empty
sysUndefinedAttrib = module
  setStateAttrib a m
  interface
