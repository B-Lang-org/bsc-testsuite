package AbstractDeriveAttrib where

a :: Attributes__
a = _

m :: Module Empty
m = module
  interface

sysAbstractDeriveAttrib :: Module Empty
sysAbstractDeriveAttrib = module
  setStateAttrib a m
  interface
